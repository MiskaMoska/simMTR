`include "params.vh"
module MTR(
    input       wire                            clk,
    input       wire                            rstn,

    input       wire        [`DW-1:0]           data_i_0_0_0,
    input       wire                            valid_i_0_0_0,
    output      wire                            ready_o_0_0_0,
    output      wire        [`DW-1:0]           data_o_0_0_0,
    output      wire                            valid_o_0_0_0,
    input       wire                            ready_i_0_0_0,

    input       wire        [`DW-1:0]           data_i_0_0_1,
    input       wire                            valid_i_0_0_1,
    output      wire                            ready_o_0_0_1,
    output      wire        [`DW-1:0]           data_o_0_0_1,
    output      wire                            valid_o_0_0_1,
    input       wire                            ready_i_0_0_1,

    input       wire        [`DW-1:0]           data_i_0_0_2,
    input       wire                            valid_i_0_0_2,
    output      wire                            ready_o_0_0_2,
    output      wire        [`DW-1:0]           data_o_0_0_2,
    output      wire                            valid_o_0_0_2,
    input       wire                            ready_i_0_0_2,

    input       wire        [`DW-1:0]           data_i_0_0_3,
    input       wire                            valid_i_0_0_3,
    output      wire                            ready_o_0_0_3,
    output      wire        [`DW-1:0]           data_o_0_0_3,
    output      wire                            valid_o_0_0_3,
    input       wire                            ready_i_0_0_3,

    input       wire        [`DW-1:0]           data_i_0_1_0,
    input       wire                            valid_i_0_1_0,
    output      wire                            ready_o_0_1_0,
    output      wire        [`DW-1:0]           data_o_0_1_0,
    output      wire                            valid_o_0_1_0,
    input       wire                            ready_i_0_1_0,

    input       wire        [`DW-1:0]           data_i_0_1_1,
    input       wire                            valid_i_0_1_1,
    output      wire                            ready_o_0_1_1,
    output      wire        [`DW-1:0]           data_o_0_1_1,
    output      wire                            valid_o_0_1_1,
    input       wire                            ready_i_0_1_1,

    input       wire        [`DW-1:0]           data_i_0_1_2,
    input       wire                            valid_i_0_1_2,
    output      wire                            ready_o_0_1_2,
    output      wire        [`DW-1:0]           data_o_0_1_2,
    output      wire                            valid_o_0_1_2,
    input       wire                            ready_i_0_1_2,

    input       wire        [`DW-1:0]           data_i_0_1_3,
    input       wire                            valid_i_0_1_3,
    output      wire                            ready_o_0_1_3,
    output      wire        [`DW-1:0]           data_o_0_1_3,
    output      wire                            valid_o_0_1_3,
    input       wire                            ready_i_0_1_3,

    input       wire        [`DW-1:0]           data_i_0_2_0,
    input       wire                            valid_i_0_2_0,
    output      wire                            ready_o_0_2_0,
    output      wire        [`DW-1:0]           data_o_0_2_0,
    output      wire                            valid_o_0_2_0,
    input       wire                            ready_i_0_2_0,

    input       wire        [`DW-1:0]           data_i_0_2_1,
    input       wire                            valid_i_0_2_1,
    output      wire                            ready_o_0_2_1,
    output      wire        [`DW-1:0]           data_o_0_2_1,
    output      wire                            valid_o_0_2_1,
    input       wire                            ready_i_0_2_1,

    input       wire        [`DW-1:0]           data_i_0_2_2,
    input       wire                            valid_i_0_2_2,
    output      wire                            ready_o_0_2_2,
    output      wire        [`DW-1:0]           data_o_0_2_2,
    output      wire                            valid_o_0_2_2,
    input       wire                            ready_i_0_2_2,

    input       wire        [`DW-1:0]           data_i_0_2_3,
    input       wire                            valid_i_0_2_3,
    output      wire                            ready_o_0_2_3,
    output      wire        [`DW-1:0]           data_o_0_2_3,
    output      wire                            valid_o_0_2_3,
    input       wire                            ready_i_0_2_3,

    input       wire        [`DW-1:0]           data_i_0_3_0,
    input       wire                            valid_i_0_3_0,
    output      wire                            ready_o_0_3_0,
    output      wire        [`DW-1:0]           data_o_0_3_0,
    output      wire                            valid_o_0_3_0,
    input       wire                            ready_i_0_3_0,

    input       wire        [`DW-1:0]           data_i_0_3_1,
    input       wire                            valid_i_0_3_1,
    output      wire                            ready_o_0_3_1,
    output      wire        [`DW-1:0]           data_o_0_3_1,
    output      wire                            valid_o_0_3_1,
    input       wire                            ready_i_0_3_1,

    input       wire        [`DW-1:0]           data_i_0_3_2,
    input       wire                            valid_i_0_3_2,
    output      wire                            ready_o_0_3_2,
    output      wire        [`DW-1:0]           data_o_0_3_2,
    output      wire                            valid_o_0_3_2,
    input       wire                            ready_i_0_3_2,

    input       wire        [`DW-1:0]           data_i_0_3_3,
    input       wire                            valid_i_0_3_3,
    output      wire                            ready_o_0_3_3,
    output      wire        [`DW-1:0]           data_o_0_3_3,
    output      wire                            valid_o_0_3_3,
    input       wire                            ready_i_0_3_3,

    input       wire        [`DW-1:0]           data_i_1_0_0,
    input       wire                            valid_i_1_0_0,
    output      wire                            ready_o_1_0_0,
    output      wire        [`DW-1:0]           data_o_1_0_0,
    output      wire                            valid_o_1_0_0,
    input       wire                            ready_i_1_0_0,

    input       wire        [`DW-1:0]           data_i_1_0_1,
    input       wire                            valid_i_1_0_1,
    output      wire                            ready_o_1_0_1,
    output      wire        [`DW-1:0]           data_o_1_0_1,
    output      wire                            valid_o_1_0_1,
    input       wire                            ready_i_1_0_1,

    input       wire        [`DW-1:0]           data_i_1_0_2,
    input       wire                            valid_i_1_0_2,
    output      wire                            ready_o_1_0_2,
    output      wire        [`DW-1:0]           data_o_1_0_2,
    output      wire                            valid_o_1_0_2,
    input       wire                            ready_i_1_0_2,

    input       wire        [`DW-1:0]           data_i_1_0_3,
    input       wire                            valid_i_1_0_3,
    output      wire                            ready_o_1_0_3,
    output      wire        [`DW-1:0]           data_o_1_0_3,
    output      wire                            valid_o_1_0_3,
    input       wire                            ready_i_1_0_3,

    input       wire        [`DW-1:0]           data_i_1_1_0,
    input       wire                            valid_i_1_1_0,
    output      wire                            ready_o_1_1_0,
    output      wire        [`DW-1:0]           data_o_1_1_0,
    output      wire                            valid_o_1_1_0,
    input       wire                            ready_i_1_1_0,

    input       wire        [`DW-1:0]           data_i_1_1_1,
    input       wire                            valid_i_1_1_1,
    output      wire                            ready_o_1_1_1,
    output      wire        [`DW-1:0]           data_o_1_1_1,
    output      wire                            valid_o_1_1_1,
    input       wire                            ready_i_1_1_1,

    input       wire        [`DW-1:0]           data_i_1_1_2,
    input       wire                            valid_i_1_1_2,
    output      wire                            ready_o_1_1_2,
    output      wire        [`DW-1:0]           data_o_1_1_2,
    output      wire                            valid_o_1_1_2,
    input       wire                            ready_i_1_1_2,

    input       wire        [`DW-1:0]           data_i_1_1_3,
    input       wire                            valid_i_1_1_3,
    output      wire                            ready_o_1_1_3,
    output      wire        [`DW-1:0]           data_o_1_1_3,
    output      wire                            valid_o_1_1_3,
    input       wire                            ready_i_1_1_3,

    input       wire        [`DW-1:0]           data_i_1_2_0,
    input       wire                            valid_i_1_2_0,
    output      wire                            ready_o_1_2_0,
    output      wire        [`DW-1:0]           data_o_1_2_0,
    output      wire                            valid_o_1_2_0,
    input       wire                            ready_i_1_2_0,

    input       wire        [`DW-1:0]           data_i_1_2_1,
    input       wire                            valid_i_1_2_1,
    output      wire                            ready_o_1_2_1,
    output      wire        [`DW-1:0]           data_o_1_2_1,
    output      wire                            valid_o_1_2_1,
    input       wire                            ready_i_1_2_1,

    input       wire        [`DW-1:0]           data_i_1_2_2,
    input       wire                            valid_i_1_2_2,
    output      wire                            ready_o_1_2_2,
    output      wire        [`DW-1:0]           data_o_1_2_2,
    output      wire                            valid_o_1_2_2,
    input       wire                            ready_i_1_2_2,

    input       wire        [`DW-1:0]           data_i_1_2_3,
    input       wire                            valid_i_1_2_3,
    output      wire                            ready_o_1_2_3,
    output      wire        [`DW-1:0]           data_o_1_2_3,
    output      wire                            valid_o_1_2_3,
    input       wire                            ready_i_1_2_3,

    input       wire        [`DW-1:0]           data_i_1_3_0,
    input       wire                            valid_i_1_3_0,
    output      wire                            ready_o_1_3_0,
    output      wire        [`DW-1:0]           data_o_1_3_0,
    output      wire                            valid_o_1_3_0,
    input       wire                            ready_i_1_3_0,

    input       wire        [`DW-1:0]           data_i_1_3_1,
    input       wire                            valid_i_1_3_1,
    output      wire                            ready_o_1_3_1,
    output      wire        [`DW-1:0]           data_o_1_3_1,
    output      wire                            valid_o_1_3_1,
    input       wire                            ready_i_1_3_1,

    input       wire        [`DW-1:0]           data_i_1_3_2,
    input       wire                            valid_i_1_3_2,
    output      wire                            ready_o_1_3_2,
    output      wire        [`DW-1:0]           data_o_1_3_2,
    output      wire                            valid_o_1_3_2,
    input       wire                            ready_i_1_3_2,

    input       wire        [`DW-1:0]           data_i_1_3_3,
    input       wire                            valid_i_1_3_3,
    output      wire                            ready_o_1_3_3,
    output      wire        [`DW-1:0]           data_o_1_3_3,
    output      wire                            valid_o_1_3_3,
    input       wire                            ready_i_1_3_3,

    input       wire        [`DW-1:0]           data_i_2_0_0,
    input       wire                            valid_i_2_0_0,
    output      wire                            ready_o_2_0_0,
    output      wire        [`DW-1:0]           data_o_2_0_0,
    output      wire                            valid_o_2_0_0,
    input       wire                            ready_i_2_0_0,

    input       wire        [`DW-1:0]           data_i_2_0_1,
    input       wire                            valid_i_2_0_1,
    output      wire                            ready_o_2_0_1,
    output      wire        [`DW-1:0]           data_o_2_0_1,
    output      wire                            valid_o_2_0_1,
    input       wire                            ready_i_2_0_1,

    input       wire        [`DW-1:0]           data_i_2_0_2,
    input       wire                            valid_i_2_0_2,
    output      wire                            ready_o_2_0_2,
    output      wire        [`DW-1:0]           data_o_2_0_2,
    output      wire                            valid_o_2_0_2,
    input       wire                            ready_i_2_0_2,

    input       wire        [`DW-1:0]           data_i_2_0_3,
    input       wire                            valid_i_2_0_3,
    output      wire                            ready_o_2_0_3,
    output      wire        [`DW-1:0]           data_o_2_0_3,
    output      wire                            valid_o_2_0_3,
    input       wire                            ready_i_2_0_3,

    input       wire        [`DW-1:0]           data_i_2_1_0,
    input       wire                            valid_i_2_1_0,
    output      wire                            ready_o_2_1_0,
    output      wire        [`DW-1:0]           data_o_2_1_0,
    output      wire                            valid_o_2_1_0,
    input       wire                            ready_i_2_1_0,

    input       wire        [`DW-1:0]           data_i_2_1_1,
    input       wire                            valid_i_2_1_1,
    output      wire                            ready_o_2_1_1,
    output      wire        [`DW-1:0]           data_o_2_1_1,
    output      wire                            valid_o_2_1_1,
    input       wire                            ready_i_2_1_1,

    input       wire        [`DW-1:0]           data_i_2_1_2,
    input       wire                            valid_i_2_1_2,
    output      wire                            ready_o_2_1_2,
    output      wire        [`DW-1:0]           data_o_2_1_2,
    output      wire                            valid_o_2_1_2,
    input       wire                            ready_i_2_1_2,

    input       wire        [`DW-1:0]           data_i_2_1_3,
    input       wire                            valid_i_2_1_3,
    output      wire                            ready_o_2_1_3,
    output      wire        [`DW-1:0]           data_o_2_1_3,
    output      wire                            valid_o_2_1_3,
    input       wire                            ready_i_2_1_3,

    input       wire        [`DW-1:0]           data_i_2_2_0,
    input       wire                            valid_i_2_2_0,
    output      wire                            ready_o_2_2_0,
    output      wire        [`DW-1:0]           data_o_2_2_0,
    output      wire                            valid_o_2_2_0,
    input       wire                            ready_i_2_2_0,

    input       wire        [`DW-1:0]           data_i_2_2_1,
    input       wire                            valid_i_2_2_1,
    output      wire                            ready_o_2_2_1,
    output      wire        [`DW-1:0]           data_o_2_2_1,
    output      wire                            valid_o_2_2_1,
    input       wire                            ready_i_2_2_1,

    input       wire        [`DW-1:0]           data_i_2_2_2,
    input       wire                            valid_i_2_2_2,
    output      wire                            ready_o_2_2_2,
    output      wire        [`DW-1:0]           data_o_2_2_2,
    output      wire                            valid_o_2_2_2,
    input       wire                            ready_i_2_2_2,

    input       wire        [`DW-1:0]           data_i_2_2_3,
    input       wire                            valid_i_2_2_3,
    output      wire                            ready_o_2_2_3,
    output      wire        [`DW-1:0]           data_o_2_2_3,
    output      wire                            valid_o_2_2_3,
    input       wire                            ready_i_2_2_3,

    input       wire        [`DW-1:0]           data_i_2_3_0,
    input       wire                            valid_i_2_3_0,
    output      wire                            ready_o_2_3_0,
    output      wire        [`DW-1:0]           data_o_2_3_0,
    output      wire                            valid_o_2_3_0,
    input       wire                            ready_i_2_3_0,

    input       wire        [`DW-1:0]           data_i_2_3_1,
    input       wire                            valid_i_2_3_1,
    output      wire                            ready_o_2_3_1,
    output      wire        [`DW-1:0]           data_o_2_3_1,
    output      wire                            valid_o_2_3_1,
    input       wire                            ready_i_2_3_1,

    input       wire        [`DW-1:0]           data_i_2_3_2,
    input       wire                            valid_i_2_3_2,
    output      wire                            ready_o_2_3_2,
    output      wire        [`DW-1:0]           data_o_2_3_2,
    output      wire                            valid_o_2_3_2,
    input       wire                            ready_i_2_3_2,

    input       wire        [`DW-1:0]           data_i_2_3_3,
    input       wire                            valid_i_2_3_3,
    output      wire                            ready_o_2_3_3,
    output      wire        [`DW-1:0]           data_o_2_3_3,
    output      wire                            valid_o_2_3_3,
    input       wire                            ready_i_2_3_3,

    input       wire        [`DW-1:0]           data_i_3_0_0,
    input       wire                            valid_i_3_0_0,
    output      wire                            ready_o_3_0_0,
    output      wire        [`DW-1:0]           data_o_3_0_0,
    output      wire                            valid_o_3_0_0,
    input       wire                            ready_i_3_0_0,

    input       wire        [`DW-1:0]           data_i_3_0_1,
    input       wire                            valid_i_3_0_1,
    output      wire                            ready_o_3_0_1,
    output      wire        [`DW-1:0]           data_o_3_0_1,
    output      wire                            valid_o_3_0_1,
    input       wire                            ready_i_3_0_1,

    input       wire        [`DW-1:0]           data_i_3_0_2,
    input       wire                            valid_i_3_0_2,
    output      wire                            ready_o_3_0_2,
    output      wire        [`DW-1:0]           data_o_3_0_2,
    output      wire                            valid_o_3_0_2,
    input       wire                            ready_i_3_0_2,

    input       wire        [`DW-1:0]           data_i_3_0_3,
    input       wire                            valid_i_3_0_3,
    output      wire                            ready_o_3_0_3,
    output      wire        [`DW-1:0]           data_o_3_0_3,
    output      wire                            valid_o_3_0_3,
    input       wire                            ready_i_3_0_3,

    input       wire        [`DW-1:0]           data_i_3_1_0,
    input       wire                            valid_i_3_1_0,
    output      wire                            ready_o_3_1_0,
    output      wire        [`DW-1:0]           data_o_3_1_0,
    output      wire                            valid_o_3_1_0,
    input       wire                            ready_i_3_1_0,

    input       wire        [`DW-1:0]           data_i_3_1_1,
    input       wire                            valid_i_3_1_1,
    output      wire                            ready_o_3_1_1,
    output      wire        [`DW-1:0]           data_o_3_1_1,
    output      wire                            valid_o_3_1_1,
    input       wire                            ready_i_3_1_1,

    input       wire        [`DW-1:0]           data_i_3_1_2,
    input       wire                            valid_i_3_1_2,
    output      wire                            ready_o_3_1_2,
    output      wire        [`DW-1:0]           data_o_3_1_2,
    output      wire                            valid_o_3_1_2,
    input       wire                            ready_i_3_1_2,

    input       wire        [`DW-1:0]           data_i_3_1_3,
    input       wire                            valid_i_3_1_3,
    output      wire                            ready_o_3_1_3,
    output      wire        [`DW-1:0]           data_o_3_1_3,
    output      wire                            valid_o_3_1_3,
    input       wire                            ready_i_3_1_3,

    input       wire        [`DW-1:0]           data_i_3_2_0,
    input       wire                            valid_i_3_2_0,
    output      wire                            ready_o_3_2_0,
    output      wire        [`DW-1:0]           data_o_3_2_0,
    output      wire                            valid_o_3_2_0,
    input       wire                            ready_i_3_2_0,

    input       wire        [`DW-1:0]           data_i_3_2_1,
    input       wire                            valid_i_3_2_1,
    output      wire                            ready_o_3_2_1,
    output      wire        [`DW-1:0]           data_o_3_2_1,
    output      wire                            valid_o_3_2_1,
    input       wire                            ready_i_3_2_1,

    input       wire        [`DW-1:0]           data_i_3_2_2,
    input       wire                            valid_i_3_2_2,
    output      wire                            ready_o_3_2_2,
    output      wire        [`DW-1:0]           data_o_3_2_2,
    output      wire                            valid_o_3_2_2,
    input       wire                            ready_i_3_2_2,

    input       wire        [`DW-1:0]           data_i_3_2_3,
    input       wire                            valid_i_3_2_3,
    output      wire                            ready_o_3_2_3,
    output      wire        [`DW-1:0]           data_o_3_2_3,
    output      wire                            valid_o_3_2_3,
    input       wire                            ready_i_3_2_3,

    input       wire        [`DW-1:0]           data_i_3_3_0,
    input       wire                            valid_i_3_3_0,
    output      wire                            ready_o_3_3_0,
    output      wire        [`DW-1:0]           data_o_3_3_0,
    output      wire                            valid_o_3_3_0,
    input       wire                            ready_i_3_3_0,

    input       wire        [`DW-1:0]           data_i_3_3_1,
    input       wire                            valid_i_3_3_1,
    output      wire                            ready_o_3_3_1,
    output      wire        [`DW-1:0]           data_o_3_3_1,
    output      wire                            valid_o_3_3_1,
    input       wire                            ready_i_3_3_1,

    input       wire        [`DW-1:0]           data_i_3_3_2,
    input       wire                            valid_i_3_3_2,
    output      wire                            ready_o_3_3_2,
    output      wire        [`DW-1:0]           data_o_3_3_2,
    output      wire                            valid_o_3_3_2,
    input       wire                            ready_i_3_3_2,

    input       wire        [`DW-1:0]           data_i_3_3_3,
    input       wire                            valid_i_3_3_3,
    output      wire                            ready_o_3_3_3,
    output      wire        [`DW-1:0]           data_o_3_3_3,
    output      wire                            valid_o_3_3_3,
    input       wire                            ready_i_3_3_3

);
wire     [`DW-1:0]       bound_itp_data_i_0;
wire                     bound_itp_valid_i_0;
wire                     bound_itp_ready_o_0;
wire     [`DW-1:0]       bound_itp_data_o_0;
wire                     bound_itp_valid_o_0;
wire                     bound_itp_ready_i_0;
wire     [`DW-1:0]       bound_trg_data_i_0;
wire                     bound_trg_valid_i_0;
wire                     bound_trg_ready_o_0;
wire     [`DW-1:0]       bound_trg_data_o_0;
wire                     bound_trg_valid_o_0;
wire                     bound_trg_ready_i_0;
wire     [`DW-1:0]       bound_itp_data_i_4;
wire                     bound_itp_valid_i_4;
wire                     bound_itp_ready_o_4;
wire     [`DW-1:0]       bound_itp_data_o_4;
wire                     bound_itp_valid_o_4;
wire                     bound_itp_ready_i_4;
wire     [`DW-1:0]       bound_trg_data_i_4;
wire                     bound_trg_valid_i_4;
wire                     bound_trg_ready_o_4;
wire     [`DW-1:0]       bound_trg_data_o_4;
wire                     bound_trg_valid_o_4;
wire                     bound_trg_ready_i_4;
wire     [`DW-1:0]       bound_itp_data_i_8;
wire                     bound_itp_valid_i_8;
wire                     bound_itp_ready_o_8;
wire     [`DW-1:0]       bound_itp_data_o_8;
wire                     bound_itp_valid_o_8;
wire                     bound_itp_ready_i_8;
wire     [`DW-1:0]       bound_trg_data_i_8;
wire                     bound_trg_valid_i_8;
wire                     bound_trg_ready_o_8;
wire     [`DW-1:0]       bound_trg_data_o_8;
wire                     bound_trg_valid_o_8;
wire                     bound_trg_ready_i_8;
wire     [`DW-1:0]       bound_itp_data_i_12;
wire                     bound_itp_valid_i_12;
wire                     bound_itp_ready_o_12;
wire     [`DW-1:0]       bound_itp_data_o_12;
wire                     bound_itp_valid_o_12;
wire                     bound_itp_ready_i_12;
wire     [`DW-1:0]       bound_trg_data_i_12;
wire                     bound_trg_valid_i_12;
wire                     bound_trg_ready_o_12;
wire     [`DW-1:0]       bound_trg_data_o_12;
wire                     bound_trg_valid_o_12;
wire                     bound_trg_ready_i_12;
wire     [`DW-1:0]       bound_itp_data_i_1;
wire                     bound_itp_valid_i_1;
wire                     bound_itp_ready_o_1;
wire     [`DW-1:0]       bound_itp_data_o_1;
wire                     bound_itp_valid_o_1;
wire                     bound_itp_ready_i_1;
wire     [`DW-1:0]       bound_trg_data_i_1;
wire                     bound_trg_valid_i_1;
wire                     bound_trg_ready_o_1;
wire     [`DW-1:0]       bound_trg_data_o_1;
wire                     bound_trg_valid_o_1;
wire                     bound_trg_ready_i_1;
wire     [`DW-1:0]       bound_itp_data_i_5;
wire                     bound_itp_valid_i_5;
wire                     bound_itp_ready_o_5;
wire     [`DW-1:0]       bound_itp_data_o_5;
wire                     bound_itp_valid_o_5;
wire                     bound_itp_ready_i_5;
wire     [`DW-1:0]       bound_trg_data_i_5;
wire                     bound_trg_valid_i_5;
wire                     bound_trg_ready_o_5;
wire     [`DW-1:0]       bound_trg_data_o_5;
wire                     bound_trg_valid_o_5;
wire                     bound_trg_ready_i_5;
wire     [`DW-1:0]       bound_itp_data_i_9;
wire                     bound_itp_valid_i_9;
wire                     bound_itp_ready_o_9;
wire     [`DW-1:0]       bound_itp_data_o_9;
wire                     bound_itp_valid_o_9;
wire                     bound_itp_ready_i_9;
wire     [`DW-1:0]       bound_trg_data_i_9;
wire                     bound_trg_valid_i_9;
wire                     bound_trg_ready_o_9;
wire     [`DW-1:0]       bound_trg_data_o_9;
wire                     bound_trg_valid_o_9;
wire                     bound_trg_ready_i_9;
wire     [`DW-1:0]       bound_itp_data_i_13;
wire                     bound_itp_valid_i_13;
wire                     bound_itp_ready_o_13;
wire     [`DW-1:0]       bound_itp_data_o_13;
wire                     bound_itp_valid_o_13;
wire                     bound_itp_ready_i_13;
wire     [`DW-1:0]       bound_trg_data_i_13;
wire                     bound_trg_valid_i_13;
wire                     bound_trg_ready_o_13;
wire     [`DW-1:0]       bound_trg_data_o_13;
wire                     bound_trg_valid_o_13;
wire                     bound_trg_ready_i_13;
wire     [`DW-1:0]       bound_itp_data_i_2;
wire                     bound_itp_valid_i_2;
wire                     bound_itp_ready_o_2;
wire     [`DW-1:0]       bound_itp_data_o_2;
wire                     bound_itp_valid_o_2;
wire                     bound_itp_ready_i_2;
wire     [`DW-1:0]       bound_trg_data_i_2;
wire                     bound_trg_valid_i_2;
wire                     bound_trg_ready_o_2;
wire     [`DW-1:0]       bound_trg_data_o_2;
wire                     bound_trg_valid_o_2;
wire                     bound_trg_ready_i_2;
wire     [`DW-1:0]       bound_itp_data_i_6;
wire                     bound_itp_valid_i_6;
wire                     bound_itp_ready_o_6;
wire     [`DW-1:0]       bound_itp_data_o_6;
wire                     bound_itp_valid_o_6;
wire                     bound_itp_ready_i_6;
wire     [`DW-1:0]       bound_trg_data_i_6;
wire                     bound_trg_valid_i_6;
wire                     bound_trg_ready_o_6;
wire     [`DW-1:0]       bound_trg_data_o_6;
wire                     bound_trg_valid_o_6;
wire                     bound_trg_ready_i_6;
wire     [`DW-1:0]       bound_itp_data_i_10;
wire                     bound_itp_valid_i_10;
wire                     bound_itp_ready_o_10;
wire     [`DW-1:0]       bound_itp_data_o_10;
wire                     bound_itp_valid_o_10;
wire                     bound_itp_ready_i_10;
wire     [`DW-1:0]       bound_trg_data_i_10;
wire                     bound_trg_valid_i_10;
wire                     bound_trg_ready_o_10;
wire     [`DW-1:0]       bound_trg_data_o_10;
wire                     bound_trg_valid_o_10;
wire                     bound_trg_ready_i_10;
wire     [`DW-1:0]       bound_itp_data_i_14;
wire                     bound_itp_valid_i_14;
wire                     bound_itp_ready_o_14;
wire     [`DW-1:0]       bound_itp_data_o_14;
wire                     bound_itp_valid_o_14;
wire                     bound_itp_ready_i_14;
wire     [`DW-1:0]       bound_trg_data_i_14;
wire                     bound_trg_valid_i_14;
wire                     bound_trg_ready_o_14;
wire     [`DW-1:0]       bound_trg_data_o_14;
wire                     bound_trg_valid_o_14;
wire                     bound_trg_ready_i_14;
wire     [`DW-1:0]       bound_itp_data_i_3;
wire                     bound_itp_valid_i_3;
wire                     bound_itp_ready_o_3;
wire     [`DW-1:0]       bound_itp_data_o_3;
wire                     bound_itp_valid_o_3;
wire                     bound_itp_ready_i_3;
wire     [`DW-1:0]       bound_trg_data_i_3;
wire                     bound_trg_valid_i_3;
wire                     bound_trg_ready_o_3;
wire     [`DW-1:0]       bound_trg_data_o_3;
wire                     bound_trg_valid_o_3;
wire                     bound_trg_ready_i_3;
wire     [`DW-1:0]       bound_itp_data_i_7;
wire                     bound_itp_valid_i_7;
wire                     bound_itp_ready_o_7;
wire     [`DW-1:0]       bound_itp_data_o_7;
wire                     bound_itp_valid_o_7;
wire                     bound_itp_ready_i_7;
wire     [`DW-1:0]       bound_trg_data_i_7;
wire                     bound_trg_valid_i_7;
wire                     bound_trg_ready_o_7;
wire     [`DW-1:0]       bound_trg_data_o_7;
wire                     bound_trg_valid_o_7;
wire                     bound_trg_ready_i_7;
wire     [`DW-1:0]       bound_itp_data_i_11;
wire                     bound_itp_valid_i_11;
wire                     bound_itp_ready_o_11;
wire     [`DW-1:0]       bound_itp_data_o_11;
wire                     bound_itp_valid_o_11;
wire                     bound_itp_ready_i_11;
wire     [`DW-1:0]       bound_trg_data_i_11;
wire                     bound_trg_valid_i_11;
wire                     bound_trg_ready_o_11;
wire     [`DW-1:0]       bound_trg_data_o_11;
wire                     bound_trg_valid_o_11;
wire                     bound_trg_ready_i_11;
wire     [`DW-1:0]       bound_itp_data_i_15;
wire                     bound_itp_valid_i_15;
wire                     bound_itp_ready_o_15;
wire     [`DW-1:0]       bound_itp_data_o_15;
wire                     bound_itp_valid_o_15;
wire                     bound_itp_ready_i_15;
wire     [`DW-1:0]       bound_trg_data_i_15;
wire                     bound_trg_valid_i_15;
wire                     bound_trg_ready_o_15;
wire     [`DW-1:0]       bound_trg_data_o_15;
wire                     bound_trg_valid_o_15;
wire                     bound_trg_ready_i_15;

InterposerNoC inoc(
    
    .clk                        (clk),
    .rstn                       (rstn),
    

    .data_i_0_0                 (bound_itp_data_i_0),
    .valid_i_0_0                (bound_itp_valid_i_0),
    .ready_o_0_0                (bound_itp_ready_o_0),
    .data_o_0_0                 (bound_itp_data_o_0),
    .valid_o_0_0                (bound_itp_valid_o_0),
    .ready_i_0_0                (bound_itp_ready_i_0),

    .data_i_0_1                 (bound_itp_data_i_4),
    .valid_i_0_1                (bound_itp_valid_i_4),
    .ready_o_0_1                (bound_itp_ready_o_4),
    .data_o_0_1                 (bound_itp_data_o_4),
    .valid_o_0_1                (bound_itp_valid_o_4),
    .ready_i_0_1                (bound_itp_ready_i_4),

    .data_i_0_2                 (bound_itp_data_i_8),
    .valid_i_0_2                (bound_itp_valid_i_8),
    .ready_o_0_2                (bound_itp_ready_o_8),
    .data_o_0_2                 (bound_itp_data_o_8),
    .valid_o_0_2                (bound_itp_valid_o_8),
    .ready_i_0_2                (bound_itp_ready_i_8),

    .data_i_0_3                 (bound_itp_data_i_12),
    .valid_i_0_3                (bound_itp_valid_i_12),
    .ready_o_0_3                (bound_itp_ready_o_12),
    .data_o_0_3                 (bound_itp_data_o_12),
    .valid_o_0_3                (bound_itp_valid_o_12),
    .ready_i_0_3                (bound_itp_ready_i_12),

    .data_i_1_0                 (bound_itp_data_i_1),
    .valid_i_1_0                (bound_itp_valid_i_1),
    .ready_o_1_0                (bound_itp_ready_o_1),
    .data_o_1_0                 (bound_itp_data_o_1),
    .valid_o_1_0                (bound_itp_valid_o_1),
    .ready_i_1_0                (bound_itp_ready_i_1),

    .data_i_1_1                 (bound_itp_data_i_5),
    .valid_i_1_1                (bound_itp_valid_i_5),
    .ready_o_1_1                (bound_itp_ready_o_5),
    .data_o_1_1                 (bound_itp_data_o_5),
    .valid_o_1_1                (bound_itp_valid_o_5),
    .ready_i_1_1                (bound_itp_ready_i_5),

    .data_i_1_2                 (bound_itp_data_i_9),
    .valid_i_1_2                (bound_itp_valid_i_9),
    .ready_o_1_2                (bound_itp_ready_o_9),
    .data_o_1_2                 (bound_itp_data_o_9),
    .valid_o_1_2                (bound_itp_valid_o_9),
    .ready_i_1_2                (bound_itp_ready_i_9),

    .data_i_1_3                 (bound_itp_data_i_13),
    .valid_i_1_3                (bound_itp_valid_i_13),
    .ready_o_1_3                (bound_itp_ready_o_13),
    .data_o_1_3                 (bound_itp_data_o_13),
    .valid_o_1_3                (bound_itp_valid_o_13),
    .ready_i_1_3                (bound_itp_ready_i_13),

    .data_i_2_0                 (bound_itp_data_i_2),
    .valid_i_2_0                (bound_itp_valid_i_2),
    .ready_o_2_0                (bound_itp_ready_o_2),
    .data_o_2_0                 (bound_itp_data_o_2),
    .valid_o_2_0                (bound_itp_valid_o_2),
    .ready_i_2_0                (bound_itp_ready_i_2),

    .data_i_2_1                 (bound_itp_data_i_6),
    .valid_i_2_1                (bound_itp_valid_i_6),
    .ready_o_2_1                (bound_itp_ready_o_6),
    .data_o_2_1                 (bound_itp_data_o_6),
    .valid_o_2_1                (bound_itp_valid_o_6),
    .ready_i_2_1                (bound_itp_ready_i_6),

    .data_i_2_2                 (bound_itp_data_i_10),
    .valid_i_2_2                (bound_itp_valid_i_10),
    .ready_o_2_2                (bound_itp_ready_o_10),
    .data_o_2_2                 (bound_itp_data_o_10),
    .valid_o_2_2                (bound_itp_valid_o_10),
    .ready_i_2_2                (bound_itp_ready_i_10),

    .data_i_2_3                 (bound_itp_data_i_14),
    .valid_i_2_3                (bound_itp_valid_i_14),
    .ready_o_2_3                (bound_itp_ready_o_14),
    .data_o_2_3                 (bound_itp_data_o_14),
    .valid_o_2_3                (bound_itp_valid_o_14),
    .ready_i_2_3                (bound_itp_ready_i_14),

    .data_i_3_0                 (bound_itp_data_i_3),
    .valid_i_3_0                (bound_itp_valid_i_3),
    .ready_o_3_0                (bound_itp_ready_o_3),
    .data_o_3_0                 (bound_itp_data_o_3),
    .valid_o_3_0                (bound_itp_valid_o_3),
    .ready_i_3_0                (bound_itp_ready_i_3),

    .data_i_3_1                 (bound_itp_data_i_7),
    .valid_i_3_1                (bound_itp_valid_i_7),
    .ready_o_3_1                (bound_itp_ready_o_7),
    .data_o_3_1                 (bound_itp_data_o_7),
    .valid_o_3_1                (bound_itp_valid_o_7),
    .ready_i_3_1                (bound_itp_ready_i_7),

    .data_i_3_2                 (bound_itp_data_i_11),
    .valid_i_3_2                (bound_itp_valid_i_11),
    .ready_o_3_2                (bound_itp_ready_o_11),
    .data_o_3_2                 (bound_itp_data_o_11),
    .valid_o_3_2                (bound_itp_valid_o_11),
    .ready_i_3_2                (bound_itp_ready_i_11),

    .data_i_3_3                 (bound_itp_data_i_15),
    .valid_i_3_3                (bound_itp_valid_i_15),
    .ready_o_3_3                (bound_itp_ready_o_15),
    .data_o_3_3                 (bound_itp_data_o_15),
    .valid_o_3_3                (bound_itp_valid_o_15),
    .ready_i_3_3                (bound_itp_ready_i_15)

);

TargetNoC tnoc0(
    
    .clk                             (clk),
    .rstn                            (rstn),
 
    .local_data_i_0_0                (data_i_0_0_0),
    .local_valid_i_0_0               (valid_i_0_0_0),
    .local_ready_o_0_0               (ready_o_0_0_0),
    .local_data_o_0_0                (data_o_0_0_0),
    .local_valid_o_0_0               (valid_o_0_0_0),
    .local_ready_i_0_0               (ready_i_0_0_0),

    .bound_data_i_0_0                (64'b0),
    .bound_valid_i_0_0               (1'b0),
    .bound_ready_o_0_0               ( ),
    .bound_data_o_0_0                ( ),
    .bound_valid_o_0_0               ( ),
    .bound_ready_i_0_0               (1'b0),
 
    .local_data_i_0_1                (data_i_0_0_1),
    .local_valid_i_0_1               (valid_i_0_0_1),
    .local_ready_o_0_1               (ready_o_0_0_1),
    .local_data_o_0_1                (data_o_0_0_1),
    .local_valid_o_0_1               (valid_o_0_0_1),
    .local_ready_i_0_1               (ready_i_0_0_1),

    .bound_data_i_0_1                (64'b0),
    .bound_valid_i_0_1               (1'b0),
    .bound_ready_o_0_1               ( ),
    .bound_data_o_0_1                ( ),
    .bound_valid_o_0_1               ( ),
    .bound_ready_i_0_1               (1'b0),
 
    .local_data_i_0_2                (data_i_0_0_2),
    .local_valid_i_0_2               (valid_i_0_0_2),
    .local_ready_o_0_2               (ready_o_0_0_2),
    .local_data_o_0_2                (data_o_0_0_2),
    .local_valid_o_0_2               (valid_o_0_0_2),
    .local_ready_i_0_2               (ready_i_0_0_2),

    .bound_data_i_0_2                (bound_trg_data_i_1),
    .bound_valid_i_0_2               (bound_trg_valid_i_1),
    .bound_ready_o_0_2               (bound_trg_ready_o_1),
    .bound_data_o_0_2                (bound_trg_data_o_1),
    .bound_valid_o_0_2               (bound_trg_valid_o_1),
    .bound_ready_i_0_2               (bound_trg_ready_i_1),
 
    .local_data_i_0_3                (data_i_0_0_3),
    .local_valid_i_0_3               (valid_i_0_0_3),
    .local_ready_o_0_3               (ready_o_0_0_3),
    .local_data_o_0_3                (data_o_0_0_3),
    .local_valid_o_0_3               (valid_o_0_0_3),
    .local_ready_i_0_3               (ready_i_0_0_3),

    .bound_data_i_0_3                (64'b0),
    .bound_valid_i_0_3               (1'b0),
    .bound_ready_o_0_3               ( ),
    .bound_data_o_0_3                ( ),
    .bound_valid_o_0_3               ( ),
    .bound_ready_i_0_3               (1'b0),
 
    .local_data_i_1_0                (data_i_0_1_0),
    .local_valid_i_1_0               (valid_i_0_1_0),
    .local_ready_o_1_0               (ready_o_0_1_0),
    .local_data_o_1_0                (data_o_0_1_0),
    .local_valid_o_1_0               (valid_o_0_1_0),
    .local_ready_i_1_0               (ready_i_0_1_0),

    .bound_data_i_1_0                (64'b0),
    .bound_valid_i_1_0               (1'b0),
    .bound_ready_o_1_0               ( ),
    .bound_data_o_1_0                ( ),
    .bound_valid_o_1_0               ( ),
    .bound_ready_i_1_0               (1'b0),
 
    .local_data_i_1_1                (data_i_0_1_1),
    .local_valid_i_1_1               (valid_i_0_1_1),
    .local_ready_o_1_1               (ready_o_0_1_1),
    .local_data_o_1_1                (data_o_0_1_1),
    .local_valid_o_1_1               (valid_o_0_1_1),
    .local_ready_i_1_1               (ready_i_0_1_1),

    .bound_data_i_1_1                (64'b0),
    .bound_valid_i_1_1               (1'b0),
    .bound_ready_o_1_1               ( ),
    .bound_data_o_1_1                ( ),
    .bound_valid_o_1_1               ( ),
    .bound_ready_i_1_1               (1'b0),
 
    .local_data_i_1_2                (data_i_0_1_2),
    .local_valid_i_1_2               (valid_i_0_1_2),
    .local_ready_o_1_2               (ready_o_0_1_2),
    .local_data_o_1_2                (data_o_0_1_2),
    .local_valid_o_1_2               (valid_o_0_1_2),
    .local_ready_i_1_2               (ready_i_0_1_2),

    .bound_data_i_1_2                (bound_trg_data_i_4),
    .bound_valid_i_1_2               (bound_trg_valid_i_4),
    .bound_ready_o_1_2               (bound_trg_ready_o_4),
    .bound_data_o_1_2                (bound_trg_data_o_4),
    .bound_valid_o_1_2               (bound_trg_valid_o_4),
    .bound_ready_i_1_2               (bound_trg_ready_i_4),
 
    .local_data_i_1_3                (data_i_0_1_3),
    .local_valid_i_1_3               (valid_i_0_1_3),
    .local_ready_o_1_3               (ready_o_0_1_3),
    .local_data_o_1_3                (data_o_0_1_3),
    .local_valid_o_1_3               (valid_o_0_1_3),
    .local_ready_i_1_3               (ready_i_0_1_3),

    .bound_data_i_1_3                (64'b0),
    .bound_valid_i_1_3               (1'b0),
    .bound_ready_o_1_3               ( ),
    .bound_data_o_1_3                ( ),
    .bound_valid_o_1_3               ( ),
    .bound_ready_i_1_3               (1'b0),
 
    .local_data_i_2_0                (data_i_0_2_0),
    .local_valid_i_2_0               (valid_i_0_2_0),
    .local_ready_o_2_0               (ready_o_0_2_0),
    .local_data_o_2_0                (data_o_0_2_0),
    .local_valid_o_2_0               (valid_o_0_2_0),
    .local_ready_i_2_0               (ready_i_0_2_0),

    .bound_data_i_2_0                (64'b0),
    .bound_valid_i_2_0               (1'b0),
    .bound_ready_o_2_0               ( ),
    .bound_data_o_2_0                ( ),
    .bound_valid_o_2_0               ( ),
    .bound_ready_i_2_0               (1'b0),
 
    .local_data_i_2_1                (data_i_0_2_1),
    .local_valid_i_2_1               (valid_i_0_2_1),
    .local_ready_o_2_1               (ready_o_0_2_1),
    .local_data_o_2_1                (data_o_0_2_1),
    .local_valid_o_2_1               (valid_o_0_2_1),
    .local_ready_i_2_1               (ready_i_0_2_1),

    .bound_data_i_2_1                (64'b0),
    .bound_valid_i_2_1               (1'b0),
    .bound_ready_o_2_1               ( ),
    .bound_data_o_2_1                ( ),
    .bound_valid_o_2_1               ( ),
    .bound_ready_i_2_1               (1'b0),
 
    .local_data_i_2_2                (data_i_0_2_2),
    .local_valid_i_2_2               (valid_i_0_2_2),
    .local_ready_o_2_2               (ready_o_0_2_2),
    .local_data_o_2_2                (data_o_0_2_2),
    .local_valid_o_2_2               (valid_o_0_2_2),
    .local_ready_i_2_2               (ready_i_0_2_2),

    .bound_data_i_2_2                (bound_trg_data_i_5),
    .bound_valid_i_2_2               (bound_trg_valid_i_5),
    .bound_ready_o_2_2               (bound_trg_ready_o_5),
    .bound_data_o_2_2                (bound_trg_data_o_5),
    .bound_valid_o_2_2               (bound_trg_valid_o_5),
    .bound_ready_i_2_2               (bound_trg_ready_i_5),
 
    .local_data_i_2_3                (data_i_0_2_3),
    .local_valid_i_2_3               (valid_i_0_2_3),
    .local_ready_o_2_3               (ready_o_0_2_3),
    .local_data_o_2_3                (data_o_0_2_3),
    .local_valid_o_2_3               (valid_o_0_2_3),
    .local_ready_i_2_3               (ready_i_0_2_3),

    .bound_data_i_2_3                (64'b0),
    .bound_valid_i_2_3               (1'b0),
    .bound_ready_o_2_3               ( ),
    .bound_data_o_2_3                ( ),
    .bound_valid_o_2_3               ( ),
    .bound_ready_i_2_3               (1'b0),
 
    .local_data_i_3_0                (data_i_0_3_0),
    .local_valid_i_3_0               (valid_i_0_3_0),
    .local_ready_o_3_0               (ready_o_0_3_0),
    .local_data_o_3_0                (data_o_0_3_0),
    .local_valid_o_3_0               (valid_o_0_3_0),
    .local_ready_i_3_0               (ready_i_0_3_0),

    .bound_data_i_3_0                (64'b0),
    .bound_valid_i_3_0               (1'b0),
    .bound_ready_o_3_0               ( ),
    .bound_data_o_3_0                ( ),
    .bound_valid_o_3_0               ( ),
    .bound_ready_i_3_0               (1'b0),
 
    .local_data_i_3_1                (data_i_0_3_1),
    .local_valid_i_3_1               (valid_i_0_3_1),
    .local_ready_o_3_1               (ready_o_0_3_1),
    .local_data_o_3_1                (data_o_0_3_1),
    .local_valid_o_3_1               (valid_o_0_3_1),
    .local_ready_i_3_1               (ready_i_0_3_1),

    .bound_data_i_3_1                (bound_trg_data_i_0),
    .bound_valid_i_3_1               (bound_trg_valid_i_0),
    .bound_ready_o_3_1               (bound_trg_ready_o_0),
    .bound_data_o_3_1                (bound_trg_data_o_0),
    .bound_valid_o_3_1               (bound_trg_valid_o_0),
    .bound_ready_i_3_1               (bound_trg_ready_i_0),
 
    .local_data_i_3_2                (data_i_0_3_2),
    .local_valid_i_3_2               (valid_i_0_3_2),
    .local_ready_o_3_2               (ready_o_0_3_2),
    .local_data_o_3_2                (data_o_0_3_2),
    .local_valid_o_3_2               (valid_o_0_3_2),
    .local_ready_i_3_2               (ready_i_0_3_2),

    .bound_data_i_3_2                (64'b0),
    .bound_valid_i_3_2               (1'b0),
    .bound_ready_o_3_2               ( ),
    .bound_data_o_3_2                ( ),
    .bound_valid_o_3_2               ( ),
    .bound_ready_i_3_2               (1'b0),
 
    .local_data_i_3_3                (data_i_0_3_3),
    .local_valid_i_3_3               (valid_i_0_3_3),
    .local_ready_o_3_3               (ready_o_0_3_3),
    .local_data_o_3_3                (data_o_0_3_3),
    .local_valid_o_3_3               (valid_o_0_3_3),
    .local_ready_i_3_3               (ready_i_0_3_3),

    .bound_data_i_3_3                (64'b0),
    .bound_valid_i_3_3               (1'b0),
    .bound_ready_o_3_3               ( ),
    .bound_data_o_3_3                ( ),
    .bound_valid_o_3_3               ( ),
    .bound_ready_i_3_3               (1'b0)

);

TargetNoC tnoc1(
    
    .clk                             (clk),
    .rstn                            (rstn),
 
    .local_data_i_0_0                (data_i_1_0_0),
    .local_valid_i_0_0               (valid_i_1_0_0),
    .local_ready_o_0_0               (ready_o_1_0_0),
    .local_data_o_0_0                (data_o_1_0_0),
    .local_valid_o_0_0               (valid_o_1_0_0),
    .local_ready_i_0_0               (ready_i_1_0_0),

    .bound_data_i_0_0                (64'b0),
    .bound_valid_i_0_0               (1'b0),
    .bound_ready_o_0_0               ( ),
    .bound_data_o_0_0                ( ),
    .bound_valid_o_0_0               ( ),
    .bound_ready_i_0_0               (1'b0),
 
    .local_data_i_0_1                (data_i_1_0_1),
    .local_valid_i_0_1               (valid_i_1_0_1),
    .local_ready_o_0_1               (ready_o_1_0_1),
    .local_data_o_0_1                (data_o_1_0_1),
    .local_valid_o_0_1               (valid_o_1_0_1),
    .local_ready_i_0_1               (ready_i_1_0_1),

    .bound_data_i_0_1                (64'b0),
    .bound_valid_i_0_1               (1'b0),
    .bound_ready_o_0_1               ( ),
    .bound_data_o_0_1                ( ),
    .bound_valid_o_0_1               ( ),
    .bound_ready_i_0_1               (1'b0),
 
    .local_data_i_0_2                (data_i_1_0_2),
    .local_valid_i_0_2               (valid_i_1_0_2),
    .local_ready_o_0_2               (ready_o_1_0_2),
    .local_data_o_0_2                (data_o_1_0_2),
    .local_valid_o_0_2               (valid_o_1_0_2),
    .local_ready_i_0_2               (ready_i_1_0_2),

    .bound_data_i_0_2                (bound_trg_data_i_3),
    .bound_valid_i_0_2               (bound_trg_valid_i_3),
    .bound_ready_o_0_2               (bound_trg_ready_o_3),
    .bound_data_o_0_2                (bound_trg_data_o_3),
    .bound_valid_o_0_2               (bound_trg_valid_o_3),
    .bound_ready_i_0_2               (bound_trg_ready_i_3),
 
    .local_data_i_0_3                (data_i_1_0_3),
    .local_valid_i_0_3               (valid_i_1_0_3),
    .local_ready_o_0_3               (ready_o_1_0_3),
    .local_data_o_0_3                (data_o_1_0_3),
    .local_valid_o_0_3               (valid_o_1_0_3),
    .local_ready_i_0_3               (ready_i_1_0_3),

    .bound_data_i_0_3                (64'b0),
    .bound_valid_i_0_3               (1'b0),
    .bound_ready_o_0_3               ( ),
    .bound_data_o_0_3                ( ),
    .bound_valid_o_0_3               ( ),
    .bound_ready_i_0_3               (1'b0),
 
    .local_data_i_1_0                (data_i_1_1_0),
    .local_valid_i_1_0               (valid_i_1_1_0),
    .local_ready_o_1_0               (ready_o_1_1_0),
    .local_data_o_1_0                (data_o_1_1_0),
    .local_valid_o_1_0               (valid_o_1_1_0),
    .local_ready_i_1_0               (ready_i_1_1_0),

    .bound_data_i_1_0                (64'b0),
    .bound_valid_i_1_0               (1'b0),
    .bound_ready_o_1_0               ( ),
    .bound_data_o_1_0                ( ),
    .bound_valid_o_1_0               ( ),
    .bound_ready_i_1_0               (1'b0),
 
    .local_data_i_1_1                (data_i_1_1_1),
    .local_valid_i_1_1               (valid_i_1_1_1),
    .local_ready_o_1_1               (ready_o_1_1_1),
    .local_data_o_1_1                (data_o_1_1_1),
    .local_valid_o_1_1               (valid_o_1_1_1),
    .local_ready_i_1_1               (ready_i_1_1_1),

    .bound_data_i_1_1                (64'b0),
    .bound_valid_i_1_1               (1'b0),
    .bound_ready_o_1_1               ( ),
    .bound_data_o_1_1                ( ),
    .bound_valid_o_1_1               ( ),
    .bound_ready_i_1_1               (1'b0),
 
    .local_data_i_1_2                (data_i_1_1_2),
    .local_valid_i_1_2               (valid_i_1_1_2),
    .local_ready_o_1_2               (ready_o_1_1_2),
    .local_data_o_1_2                (data_o_1_1_2),
    .local_valid_o_1_2               (valid_o_1_1_2),
    .local_ready_i_1_2               (ready_i_1_1_2),

    .bound_data_i_1_2                (bound_trg_data_i_6),
    .bound_valid_i_1_2               (bound_trg_valid_i_6),
    .bound_ready_o_1_2               (bound_trg_ready_o_6),
    .bound_data_o_1_2                (bound_trg_data_o_6),
    .bound_valid_o_1_2               (bound_trg_valid_o_6),
    .bound_ready_i_1_2               (bound_trg_ready_i_6),
 
    .local_data_i_1_3                (data_i_1_1_3),
    .local_valid_i_1_3               (valid_i_1_1_3),
    .local_ready_o_1_3               (ready_o_1_1_3),
    .local_data_o_1_3                (data_o_1_1_3),
    .local_valid_o_1_3               (valid_o_1_1_3),
    .local_ready_i_1_3               (ready_i_1_1_3),

    .bound_data_i_1_3                (64'b0),
    .bound_valid_i_1_3               (1'b0),
    .bound_ready_o_1_3               ( ),
    .bound_data_o_1_3                ( ),
    .bound_valid_o_1_3               ( ),
    .bound_ready_i_1_3               (1'b0),
 
    .local_data_i_2_0                (data_i_1_2_0),
    .local_valid_i_2_0               (valid_i_1_2_0),
    .local_ready_o_2_0               (ready_o_1_2_0),
    .local_data_o_2_0                (data_o_1_2_0),
    .local_valid_o_2_0               (valid_o_1_2_0),
    .local_ready_i_2_0               (ready_i_1_2_0),

    .bound_data_i_2_0                (64'b0),
    .bound_valid_i_2_0               (1'b0),
    .bound_ready_o_2_0               ( ),
    .bound_data_o_2_0                ( ),
    .bound_valid_o_2_0               ( ),
    .bound_ready_i_2_0               (1'b0),
 
    .local_data_i_2_1                (data_i_1_2_1),
    .local_valid_i_2_1               (valid_i_1_2_1),
    .local_ready_o_2_1               (ready_o_1_2_1),
    .local_data_o_2_1                (data_o_1_2_1),
    .local_valid_o_2_1               (valid_o_1_2_1),
    .local_ready_i_2_1               (ready_i_1_2_1),

    .bound_data_i_2_1                (64'b0),
    .bound_valid_i_2_1               (1'b0),
    .bound_ready_o_2_1               ( ),
    .bound_data_o_2_1                ( ),
    .bound_valid_o_2_1               ( ),
    .bound_ready_i_2_1               (1'b0),
 
    .local_data_i_2_2                (data_i_1_2_2),
    .local_valid_i_2_2               (valid_i_1_2_2),
    .local_ready_o_2_2               (ready_o_1_2_2),
    .local_data_o_2_2                (data_o_1_2_2),
    .local_valid_o_2_2               (valid_o_1_2_2),
    .local_ready_i_2_2               (ready_i_1_2_2),

    .bound_data_i_2_2                (bound_trg_data_i_7),
    .bound_valid_i_2_2               (bound_trg_valid_i_7),
    .bound_ready_o_2_2               (bound_trg_ready_o_7),
    .bound_data_o_2_2                (bound_trg_data_o_7),
    .bound_valid_o_2_2               (bound_trg_valid_o_7),
    .bound_ready_i_2_2               (bound_trg_ready_i_7),
 
    .local_data_i_2_3                (data_i_1_2_3),
    .local_valid_i_2_3               (valid_i_1_2_3),
    .local_ready_o_2_3               (ready_o_1_2_3),
    .local_data_o_2_3                (data_o_1_2_3),
    .local_valid_o_2_3               (valid_o_1_2_3),
    .local_ready_i_2_3               (ready_i_1_2_3),

    .bound_data_i_2_3                (64'b0),
    .bound_valid_i_2_3               (1'b0),
    .bound_ready_o_2_3               ( ),
    .bound_data_o_2_3                ( ),
    .bound_valid_o_2_3               ( ),
    .bound_ready_i_2_3               (1'b0),
 
    .local_data_i_3_0                (data_i_1_3_0),
    .local_valid_i_3_0               (valid_i_1_3_0),
    .local_ready_o_3_0               (ready_o_1_3_0),
    .local_data_o_3_0                (data_o_1_3_0),
    .local_valid_o_3_0               (valid_o_1_3_0),
    .local_ready_i_3_0               (ready_i_1_3_0),

    .bound_data_i_3_0                (64'b0),
    .bound_valid_i_3_0               (1'b0),
    .bound_ready_o_3_0               ( ),
    .bound_data_o_3_0                ( ),
    .bound_valid_o_3_0               ( ),
    .bound_ready_i_3_0               (1'b0),
 
    .local_data_i_3_1                (data_i_1_3_1),
    .local_valid_i_3_1               (valid_i_1_3_1),
    .local_ready_o_3_1               (ready_o_1_3_1),
    .local_data_o_3_1                (data_o_1_3_1),
    .local_valid_o_3_1               (valid_o_1_3_1),
    .local_ready_i_3_1               (ready_i_1_3_1),

    .bound_data_i_3_1                (bound_trg_data_i_2),
    .bound_valid_i_3_1               (bound_trg_valid_i_2),
    .bound_ready_o_3_1               (bound_trg_ready_o_2),
    .bound_data_o_3_1                (bound_trg_data_o_2),
    .bound_valid_o_3_1               (bound_trg_valid_o_2),
    .bound_ready_i_3_1               (bound_trg_ready_i_2),
 
    .local_data_i_3_2                (data_i_1_3_2),
    .local_valid_i_3_2               (valid_i_1_3_2),
    .local_ready_o_3_2               (ready_o_1_3_2),
    .local_data_o_3_2                (data_o_1_3_2),
    .local_valid_o_3_2               (valid_o_1_3_2),
    .local_ready_i_3_2               (ready_i_1_3_2),

    .bound_data_i_3_2                (64'b0),
    .bound_valid_i_3_2               (1'b0),
    .bound_ready_o_3_2               ( ),
    .bound_data_o_3_2                ( ),
    .bound_valid_o_3_2               ( ),
    .bound_ready_i_3_2               (1'b0),
 
    .local_data_i_3_3                (data_i_1_3_3),
    .local_valid_i_3_3               (valid_i_1_3_3),
    .local_ready_o_3_3               (ready_o_1_3_3),
    .local_data_o_3_3                (data_o_1_3_3),
    .local_valid_o_3_3               (valid_o_1_3_3),
    .local_ready_i_3_3               (ready_i_1_3_3),

    .bound_data_i_3_3                (64'b0),
    .bound_valid_i_3_3               (1'b0),
    .bound_ready_o_3_3               ( ),
    .bound_data_o_3_3                ( ),
    .bound_valid_o_3_3               ( ),
    .bound_ready_i_3_3               (1'b0)

);

TargetNoC tnoc2(
    
    .clk                             (clk),
    .rstn                            (rstn),
 
    .local_data_i_0_0                (data_i_2_0_0),
    .local_valid_i_0_0               (valid_i_2_0_0),
    .local_ready_o_0_0               (ready_o_2_0_0),
    .local_data_o_0_0                (data_o_2_0_0),
    .local_valid_o_0_0               (valid_o_2_0_0),
    .local_ready_i_0_0               (ready_i_2_0_0),

    .bound_data_i_0_0                (64'b0),
    .bound_valid_i_0_0               (1'b0),
    .bound_ready_o_0_0               ( ),
    .bound_data_o_0_0                ( ),
    .bound_valid_o_0_0               ( ),
    .bound_ready_i_0_0               (1'b0),
 
    .local_data_i_0_1                (data_i_2_0_1),
    .local_valid_i_0_1               (valid_i_2_0_1),
    .local_ready_o_0_1               (ready_o_2_0_1),
    .local_data_o_0_1                (data_o_2_0_1),
    .local_valid_o_0_1               (valid_o_2_0_1),
    .local_ready_i_0_1               (ready_i_2_0_1),

    .bound_data_i_0_1                (64'b0),
    .bound_valid_i_0_1               (1'b0),
    .bound_ready_o_0_1               ( ),
    .bound_data_o_0_1                ( ),
    .bound_valid_o_0_1               ( ),
    .bound_ready_i_0_1               (1'b0),
 
    .local_data_i_0_2                (data_i_2_0_2),
    .local_valid_i_0_2               (valid_i_2_0_2),
    .local_ready_o_0_2               (ready_o_2_0_2),
    .local_data_o_0_2                (data_o_2_0_2),
    .local_valid_o_0_2               (valid_o_2_0_2),
    .local_ready_i_0_2               (ready_i_2_0_2),

    .bound_data_i_0_2                (bound_trg_data_i_9),
    .bound_valid_i_0_2               (bound_trg_valid_i_9),
    .bound_ready_o_0_2               (bound_trg_ready_o_9),
    .bound_data_o_0_2                (bound_trg_data_o_9),
    .bound_valid_o_0_2               (bound_trg_valid_o_9),
    .bound_ready_i_0_2               (bound_trg_ready_i_9),
 
    .local_data_i_0_3                (data_i_2_0_3),
    .local_valid_i_0_3               (valid_i_2_0_3),
    .local_ready_o_0_3               (ready_o_2_0_3),
    .local_data_o_0_3                (data_o_2_0_3),
    .local_valid_o_0_3               (valid_o_2_0_3),
    .local_ready_i_0_3               (ready_i_2_0_3),

    .bound_data_i_0_3                (64'b0),
    .bound_valid_i_0_3               (1'b0),
    .bound_ready_o_0_3               ( ),
    .bound_data_o_0_3                ( ),
    .bound_valid_o_0_3               ( ),
    .bound_ready_i_0_3               (1'b0),
 
    .local_data_i_1_0                (data_i_2_1_0),
    .local_valid_i_1_0               (valid_i_2_1_0),
    .local_ready_o_1_0               (ready_o_2_1_0),
    .local_data_o_1_0                (data_o_2_1_0),
    .local_valid_o_1_0               (valid_o_2_1_0),
    .local_ready_i_1_0               (ready_i_2_1_0),

    .bound_data_i_1_0                (64'b0),
    .bound_valid_i_1_0               (1'b0),
    .bound_ready_o_1_0               ( ),
    .bound_data_o_1_0                ( ),
    .bound_valid_o_1_0               ( ),
    .bound_ready_i_1_0               (1'b0),
 
    .local_data_i_1_1                (data_i_2_1_1),
    .local_valid_i_1_1               (valid_i_2_1_1),
    .local_ready_o_1_1               (ready_o_2_1_1),
    .local_data_o_1_1                (data_o_2_1_1),
    .local_valid_o_1_1               (valid_o_2_1_1),
    .local_ready_i_1_1               (ready_i_2_1_1),

    .bound_data_i_1_1                (64'b0),
    .bound_valid_i_1_1               (1'b0),
    .bound_ready_o_1_1               ( ),
    .bound_data_o_1_1                ( ),
    .bound_valid_o_1_1               ( ),
    .bound_ready_i_1_1               (1'b0),
 
    .local_data_i_1_2                (data_i_2_1_2),
    .local_valid_i_1_2               (valid_i_2_1_2),
    .local_ready_o_1_2               (ready_o_2_1_2),
    .local_data_o_1_2                (data_o_2_1_2),
    .local_valid_o_1_2               (valid_o_2_1_2),
    .local_ready_i_1_2               (ready_i_2_1_2),

    .bound_data_i_1_2                (bound_trg_data_i_12),
    .bound_valid_i_1_2               (bound_trg_valid_i_12),
    .bound_ready_o_1_2               (bound_trg_ready_o_12),
    .bound_data_o_1_2                (bound_trg_data_o_12),
    .bound_valid_o_1_2               (bound_trg_valid_o_12),
    .bound_ready_i_1_2               (bound_trg_ready_i_12),
 
    .local_data_i_1_3                (data_i_2_1_3),
    .local_valid_i_1_3               (valid_i_2_1_3),
    .local_ready_o_1_3               (ready_o_2_1_3),
    .local_data_o_1_3                (data_o_2_1_3),
    .local_valid_o_1_3               (valid_o_2_1_3),
    .local_ready_i_1_3               (ready_i_2_1_3),

    .bound_data_i_1_3                (64'b0),
    .bound_valid_i_1_3               (1'b0),
    .bound_ready_o_1_3               ( ),
    .bound_data_o_1_3                ( ),
    .bound_valid_o_1_3               ( ),
    .bound_ready_i_1_3               (1'b0),
 
    .local_data_i_2_0                (data_i_2_2_0),
    .local_valid_i_2_0               (valid_i_2_2_0),
    .local_ready_o_2_0               (ready_o_2_2_0),
    .local_data_o_2_0                (data_o_2_2_0),
    .local_valid_o_2_0               (valid_o_2_2_0),
    .local_ready_i_2_0               (ready_i_2_2_0),

    .bound_data_i_2_0                (64'b0),
    .bound_valid_i_2_0               (1'b0),
    .bound_ready_o_2_0               ( ),
    .bound_data_o_2_0                ( ),
    .bound_valid_o_2_0               ( ),
    .bound_ready_i_2_0               (1'b0),
 
    .local_data_i_2_1                (data_i_2_2_1),
    .local_valid_i_2_1               (valid_i_2_2_1),
    .local_ready_o_2_1               (ready_o_2_2_1),
    .local_data_o_2_1                (data_o_2_2_1),
    .local_valid_o_2_1               (valid_o_2_2_1),
    .local_ready_i_2_1               (ready_i_2_2_1),

    .bound_data_i_2_1                (64'b0),
    .bound_valid_i_2_1               (1'b0),
    .bound_ready_o_2_1               ( ),
    .bound_data_o_2_1                ( ),
    .bound_valid_o_2_1               ( ),
    .bound_ready_i_2_1               (1'b0),
 
    .local_data_i_2_2                (data_i_2_2_2),
    .local_valid_i_2_2               (valid_i_2_2_2),
    .local_ready_o_2_2               (ready_o_2_2_2),
    .local_data_o_2_2                (data_o_2_2_2),
    .local_valid_o_2_2               (valid_o_2_2_2),
    .local_ready_i_2_2               (ready_i_2_2_2),

    .bound_data_i_2_2                (bound_trg_data_i_13),
    .bound_valid_i_2_2               (bound_trg_valid_i_13),
    .bound_ready_o_2_2               (bound_trg_ready_o_13),
    .bound_data_o_2_2                (bound_trg_data_o_13),
    .bound_valid_o_2_2               (bound_trg_valid_o_13),
    .bound_ready_i_2_2               (bound_trg_ready_i_13),
 
    .local_data_i_2_3                (data_i_2_2_3),
    .local_valid_i_2_3               (valid_i_2_2_3),
    .local_ready_o_2_3               (ready_o_2_2_3),
    .local_data_o_2_3                (data_o_2_2_3),
    .local_valid_o_2_3               (valid_o_2_2_3),
    .local_ready_i_2_3               (ready_i_2_2_3),

    .bound_data_i_2_3                (64'b0),
    .bound_valid_i_2_3               (1'b0),
    .bound_ready_o_2_3               ( ),
    .bound_data_o_2_3                ( ),
    .bound_valid_o_2_3               ( ),
    .bound_ready_i_2_3               (1'b0),
 
    .local_data_i_3_0                (data_i_2_3_0),
    .local_valid_i_3_0               (valid_i_2_3_0),
    .local_ready_o_3_0               (ready_o_2_3_0),
    .local_data_o_3_0                (data_o_2_3_0),
    .local_valid_o_3_0               (valid_o_2_3_0),
    .local_ready_i_3_0               (ready_i_2_3_0),

    .bound_data_i_3_0                (64'b0),
    .bound_valid_i_3_0               (1'b0),
    .bound_ready_o_3_0               ( ),
    .bound_data_o_3_0                ( ),
    .bound_valid_o_3_0               ( ),
    .bound_ready_i_3_0               (1'b0),
 
    .local_data_i_3_1                (data_i_2_3_1),
    .local_valid_i_3_1               (valid_i_2_3_1),
    .local_ready_o_3_1               (ready_o_2_3_1),
    .local_data_o_3_1                (data_o_2_3_1),
    .local_valid_o_3_1               (valid_o_2_3_1),
    .local_ready_i_3_1               (ready_i_2_3_1),

    .bound_data_i_3_1                (bound_trg_data_i_8),
    .bound_valid_i_3_1               (bound_trg_valid_i_8),
    .bound_ready_o_3_1               (bound_trg_ready_o_8),
    .bound_data_o_3_1                (bound_trg_data_o_8),
    .bound_valid_o_3_1               (bound_trg_valid_o_8),
    .bound_ready_i_3_1               (bound_trg_ready_i_8),
 
    .local_data_i_3_2                (data_i_2_3_2),
    .local_valid_i_3_2               (valid_i_2_3_2),
    .local_ready_o_3_2               (ready_o_2_3_2),
    .local_data_o_3_2                (data_o_2_3_2),
    .local_valid_o_3_2               (valid_o_2_3_2),
    .local_ready_i_3_2               (ready_i_2_3_2),

    .bound_data_i_3_2                (64'b0),
    .bound_valid_i_3_2               (1'b0),
    .bound_ready_o_3_2               ( ),
    .bound_data_o_3_2                ( ),
    .bound_valid_o_3_2               ( ),
    .bound_ready_i_3_2               (1'b0),
 
    .local_data_i_3_3                (data_i_2_3_3),
    .local_valid_i_3_3               (valid_i_2_3_3),
    .local_ready_o_3_3               (ready_o_2_3_3),
    .local_data_o_3_3                (data_o_2_3_3),
    .local_valid_o_3_3               (valid_o_2_3_3),
    .local_ready_i_3_3               (ready_i_2_3_3),

    .bound_data_i_3_3                (64'b0),
    .bound_valid_i_3_3               (1'b0),
    .bound_ready_o_3_3               ( ),
    .bound_data_o_3_3                ( ),
    .bound_valid_o_3_3               ( ),
    .bound_ready_i_3_3               (1'b0)

);

TargetNoC tnoc3(
    
    .clk                             (clk),
    .rstn                            (rstn),
 
    .local_data_i_0_0                (data_i_3_0_0),
    .local_valid_i_0_0               (valid_i_3_0_0),
    .local_ready_o_0_0               (ready_o_3_0_0),
    .local_data_o_0_0                (data_o_3_0_0),
    .local_valid_o_0_0               (valid_o_3_0_0),
    .local_ready_i_0_0               (ready_i_3_0_0),

    .bound_data_i_0_0                (64'b0),
    .bound_valid_i_0_0               (1'b0),
    .bound_ready_o_0_0               ( ),
    .bound_data_o_0_0                ( ),
    .bound_valid_o_0_0               ( ),
    .bound_ready_i_0_0               (1'b0),
 
    .local_data_i_0_1                (data_i_3_0_1),
    .local_valid_i_0_1               (valid_i_3_0_1),
    .local_ready_o_0_1               (ready_o_3_0_1),
    .local_data_o_0_1                (data_o_3_0_1),
    .local_valid_o_0_1               (valid_o_3_0_1),
    .local_ready_i_0_1               (ready_i_3_0_1),

    .bound_data_i_0_1                (64'b0),
    .bound_valid_i_0_1               (1'b0),
    .bound_ready_o_0_1               ( ),
    .bound_data_o_0_1                ( ),
    .bound_valid_o_0_1               ( ),
    .bound_ready_i_0_1               (1'b0),
 
    .local_data_i_0_2                (data_i_3_0_2),
    .local_valid_i_0_2               (valid_i_3_0_2),
    .local_ready_o_0_2               (ready_o_3_0_2),
    .local_data_o_0_2                (data_o_3_0_2),
    .local_valid_o_0_2               (valid_o_3_0_2),
    .local_ready_i_0_2               (ready_i_3_0_2),

    .bound_data_i_0_2                (bound_trg_data_i_11),
    .bound_valid_i_0_2               (bound_trg_valid_i_11),
    .bound_ready_o_0_2               (bound_trg_ready_o_11),
    .bound_data_o_0_2                (bound_trg_data_o_11),
    .bound_valid_o_0_2               (bound_trg_valid_o_11),
    .bound_ready_i_0_2               (bound_trg_ready_i_11),
 
    .local_data_i_0_3                (data_i_3_0_3),
    .local_valid_i_0_3               (valid_i_3_0_3),
    .local_ready_o_0_3               (ready_o_3_0_3),
    .local_data_o_0_3                (data_o_3_0_3),
    .local_valid_o_0_3               (valid_o_3_0_3),
    .local_ready_i_0_3               (ready_i_3_0_3),

    .bound_data_i_0_3                (64'b0),
    .bound_valid_i_0_3               (1'b0),
    .bound_ready_o_0_3               ( ),
    .bound_data_o_0_3                ( ),
    .bound_valid_o_0_3               ( ),
    .bound_ready_i_0_3               (1'b0),
 
    .local_data_i_1_0                (data_i_3_1_0),
    .local_valid_i_1_0               (valid_i_3_1_0),
    .local_ready_o_1_0               (ready_o_3_1_0),
    .local_data_o_1_0                (data_o_3_1_0),
    .local_valid_o_1_0               (valid_o_3_1_0),
    .local_ready_i_1_0               (ready_i_3_1_0),

    .bound_data_i_1_0                (64'b0),
    .bound_valid_i_1_0               (1'b0),
    .bound_ready_o_1_0               ( ),
    .bound_data_o_1_0                ( ),
    .bound_valid_o_1_0               ( ),
    .bound_ready_i_1_0               (1'b0),
 
    .local_data_i_1_1                (data_i_3_1_1),
    .local_valid_i_1_1               (valid_i_3_1_1),
    .local_ready_o_1_1               (ready_o_3_1_1),
    .local_data_o_1_1                (data_o_3_1_1),
    .local_valid_o_1_1               (valid_o_3_1_1),
    .local_ready_i_1_1               (ready_i_3_1_1),

    .bound_data_i_1_1                (64'b0),
    .bound_valid_i_1_1               (1'b0),
    .bound_ready_o_1_1               ( ),
    .bound_data_o_1_1                ( ),
    .bound_valid_o_1_1               ( ),
    .bound_ready_i_1_1               (1'b0),
 
    .local_data_i_1_2                (data_i_3_1_2),
    .local_valid_i_1_2               (valid_i_3_1_2),
    .local_ready_o_1_2               (ready_o_3_1_2),
    .local_data_o_1_2                (data_o_3_1_2),
    .local_valid_o_1_2               (valid_o_3_1_2),
    .local_ready_i_1_2               (ready_i_3_1_2),

    .bound_data_i_1_2                (bound_trg_data_i_14),
    .bound_valid_i_1_2               (bound_trg_valid_i_14),
    .bound_ready_o_1_2               (bound_trg_ready_o_14),
    .bound_data_o_1_2                (bound_trg_data_o_14),
    .bound_valid_o_1_2               (bound_trg_valid_o_14),
    .bound_ready_i_1_2               (bound_trg_ready_i_14),
 
    .local_data_i_1_3                (data_i_3_1_3),
    .local_valid_i_1_3               (valid_i_3_1_3),
    .local_ready_o_1_3               (ready_o_3_1_3),
    .local_data_o_1_3                (data_o_3_1_3),
    .local_valid_o_1_3               (valid_o_3_1_3),
    .local_ready_i_1_3               (ready_i_3_1_3),

    .bound_data_i_1_3                (64'b0),
    .bound_valid_i_1_3               (1'b0),
    .bound_ready_o_1_3               ( ),
    .bound_data_o_1_3                ( ),
    .bound_valid_o_1_3               ( ),
    .bound_ready_i_1_3               (1'b0),
 
    .local_data_i_2_0                (data_i_3_2_0),
    .local_valid_i_2_0               (valid_i_3_2_0),
    .local_ready_o_2_0               (ready_o_3_2_0),
    .local_data_o_2_0                (data_o_3_2_0),
    .local_valid_o_2_0               (valid_o_3_2_0),
    .local_ready_i_2_0               (ready_i_3_2_0),

    .bound_data_i_2_0                (64'b0),
    .bound_valid_i_2_0               (1'b0),
    .bound_ready_o_2_0               ( ),
    .bound_data_o_2_0                ( ),
    .bound_valid_o_2_0               ( ),
    .bound_ready_i_2_0               (1'b0),
 
    .local_data_i_2_1                (data_i_3_2_1),
    .local_valid_i_2_1               (valid_i_3_2_1),
    .local_ready_o_2_1               (ready_o_3_2_1),
    .local_data_o_2_1                (data_o_3_2_1),
    .local_valid_o_2_1               (valid_o_3_2_1),
    .local_ready_i_2_1               (ready_i_3_2_1),

    .bound_data_i_2_1                (64'b0),
    .bound_valid_i_2_1               (1'b0),
    .bound_ready_o_2_1               ( ),
    .bound_data_o_2_1                ( ),
    .bound_valid_o_2_1               ( ),
    .bound_ready_i_2_1               (1'b0),
 
    .local_data_i_2_2                (data_i_3_2_2),
    .local_valid_i_2_2               (valid_i_3_2_2),
    .local_ready_o_2_2               (ready_o_3_2_2),
    .local_data_o_2_2                (data_o_3_2_2),
    .local_valid_o_2_2               (valid_o_3_2_2),
    .local_ready_i_2_2               (ready_i_3_2_2),

    .bound_data_i_2_2                (bound_trg_data_i_15),
    .bound_valid_i_2_2               (bound_trg_valid_i_15),
    .bound_ready_o_2_2               (bound_trg_ready_o_15),
    .bound_data_o_2_2                (bound_trg_data_o_15),
    .bound_valid_o_2_2               (bound_trg_valid_o_15),
    .bound_ready_i_2_2               (bound_trg_ready_i_15),
 
    .local_data_i_2_3                (data_i_3_2_3),
    .local_valid_i_2_3               (valid_i_3_2_3),
    .local_ready_o_2_3               (ready_o_3_2_3),
    .local_data_o_2_3                (data_o_3_2_3),
    .local_valid_o_2_3               (valid_o_3_2_3),
    .local_ready_i_2_3               (ready_i_3_2_3),

    .bound_data_i_2_3                (64'b0),
    .bound_valid_i_2_3               (1'b0),
    .bound_ready_o_2_3               ( ),
    .bound_data_o_2_3                ( ),
    .bound_valid_o_2_3               ( ),
    .bound_ready_i_2_3               (1'b0),
 
    .local_data_i_3_0                (data_i_3_3_0),
    .local_valid_i_3_0               (valid_i_3_3_0),
    .local_ready_o_3_0               (ready_o_3_3_0),
    .local_data_o_3_0                (data_o_3_3_0),
    .local_valid_o_3_0               (valid_o_3_3_0),
    .local_ready_i_3_0               (ready_i_3_3_0),

    .bound_data_i_3_0                (64'b0),
    .bound_valid_i_3_0               (1'b0),
    .bound_ready_o_3_0               ( ),
    .bound_data_o_3_0                ( ),
    .bound_valid_o_3_0               ( ),
    .bound_ready_i_3_0               (1'b0),
 
    .local_data_i_3_1                (data_i_3_3_1),
    .local_valid_i_3_1               (valid_i_3_3_1),
    .local_ready_o_3_1               (ready_o_3_3_1),
    .local_data_o_3_1                (data_o_3_3_1),
    .local_valid_o_3_1               (valid_o_3_3_1),
    .local_ready_i_3_1               (ready_i_3_3_1),

    .bound_data_i_3_1                (bound_trg_data_i_10),
    .bound_valid_i_3_1               (bound_trg_valid_i_10),
    .bound_ready_o_3_1               (bound_trg_ready_o_10),
    .bound_data_o_3_1                (bound_trg_data_o_10),
    .bound_valid_o_3_1               (bound_trg_valid_o_10),
    .bound_ready_i_3_1               (bound_trg_ready_i_10),
 
    .local_data_i_3_2                (data_i_3_3_2),
    .local_valid_i_3_2               (valid_i_3_3_2),
    .local_ready_o_3_2               (ready_o_3_3_2),
    .local_data_o_3_2                (data_o_3_3_2),
    .local_valid_o_3_2               (valid_o_3_3_2),
    .local_ready_i_3_2               (ready_i_3_3_2),

    .bound_data_i_3_2                (64'b0),
    .bound_valid_i_3_2               (1'b0),
    .bound_ready_o_3_2               ( ),
    .bound_data_o_3_2                ( ),
    .bound_valid_o_3_2               ( ),
    .bound_ready_i_3_2               (1'b0),
 
    .local_data_i_3_3                (data_i_3_3_3),
    .local_valid_i_3_3               (valid_i_3_3_3),
    .local_ready_o_3_3               (ready_o_3_3_3),
    .local_data_o_3_3                (data_o_3_3_3),
    .local_valid_o_3_3               (valid_o_3_3_3),
    .local_ready_i_3_3               (ready_i_3_3_3),

    .bound_data_i_3_3                (64'b0),
    .bound_valid_i_3_3               (1'b0),
    .bound_ready_o_3_3               ( ),
    .bound_data_o_3_3                ( ),
    .bound_valid_o_3_3               ( ),
    .bound_ready_i_3_3               (1'b0)

);

bound_link bl0(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_0),
    .trg_valid_i               (bound_trg_valid_o_0),
    .trg_ready_o               (bound_trg_ready_i_0),
    .trg_data_o                (bound_trg_data_i_0),
    .trg_valid_o               (bound_trg_valid_i_0),
    .trg_ready_i               (bound_trg_ready_o_0),
    .itp_data_i                (bound_itp_data_o_0),
    .itp_valid_i               (bound_itp_valid_o_0),
    .itp_ready_o               (bound_itp_ready_i_0),
    .itp_data_o                (bound_itp_data_i_0),
    .itp_valid_o               (bound_itp_valid_i_0),
    .itp_ready_i               (bound_itp_ready_o_0)
);

bound_link bl1(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_1),
    .trg_valid_i               (bound_trg_valid_o_1),
    .trg_ready_o               (bound_trg_ready_i_1),
    .trg_data_o                (bound_trg_data_i_1),
    .trg_valid_o               (bound_trg_valid_i_1),
    .trg_ready_i               (bound_trg_ready_o_1),
    .itp_data_i                (bound_itp_data_o_1),
    .itp_valid_i               (bound_itp_valid_o_1),
    .itp_ready_o               (bound_itp_ready_i_1),
    .itp_data_o                (bound_itp_data_i_1),
    .itp_valid_o               (bound_itp_valid_i_1),
    .itp_ready_i               (bound_itp_ready_o_1)
);

bound_link bl2(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_2),
    .trg_valid_i               (bound_trg_valid_o_2),
    .trg_ready_o               (bound_trg_ready_i_2),
    .trg_data_o                (bound_trg_data_i_2),
    .trg_valid_o               (bound_trg_valid_i_2),
    .trg_ready_i               (bound_trg_ready_o_2),
    .itp_data_i                (bound_itp_data_o_2),
    .itp_valid_i               (bound_itp_valid_o_2),
    .itp_ready_o               (bound_itp_ready_i_2),
    .itp_data_o                (bound_itp_data_i_2),
    .itp_valid_o               (bound_itp_valid_i_2),
    .itp_ready_i               (bound_itp_ready_o_2)
);

bound_link bl3(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_3),
    .trg_valid_i               (bound_trg_valid_o_3),
    .trg_ready_o               (bound_trg_ready_i_3),
    .trg_data_o                (bound_trg_data_i_3),
    .trg_valid_o               (bound_trg_valid_i_3),
    .trg_ready_i               (bound_trg_ready_o_3),
    .itp_data_i                (bound_itp_data_o_3),
    .itp_valid_i               (bound_itp_valid_o_3),
    .itp_ready_o               (bound_itp_ready_i_3),
    .itp_data_o                (bound_itp_data_i_3),
    .itp_valid_o               (bound_itp_valid_i_3),
    .itp_ready_i               (bound_itp_ready_o_3)
);

bound_link bl4(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_4),
    .trg_valid_i               (bound_trg_valid_o_4),
    .trg_ready_o               (bound_trg_ready_i_4),
    .trg_data_o                (bound_trg_data_i_4),
    .trg_valid_o               (bound_trg_valid_i_4),
    .trg_ready_i               (bound_trg_ready_o_4),
    .itp_data_i                (bound_itp_data_o_4),
    .itp_valid_i               (bound_itp_valid_o_4),
    .itp_ready_o               (bound_itp_ready_i_4),
    .itp_data_o                (bound_itp_data_i_4),
    .itp_valid_o               (bound_itp_valid_i_4),
    .itp_ready_i               (bound_itp_ready_o_4)
);

bound_link bl5(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_5),
    .trg_valid_i               (bound_trg_valid_o_5),
    .trg_ready_o               (bound_trg_ready_i_5),
    .trg_data_o                (bound_trg_data_i_5),
    .trg_valid_o               (bound_trg_valid_i_5),
    .trg_ready_i               (bound_trg_ready_o_5),
    .itp_data_i                (bound_itp_data_o_5),
    .itp_valid_i               (bound_itp_valid_o_5),
    .itp_ready_o               (bound_itp_ready_i_5),
    .itp_data_o                (bound_itp_data_i_5),
    .itp_valid_o               (bound_itp_valid_i_5),
    .itp_ready_i               (bound_itp_ready_o_5)
);

bound_link bl6(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_6),
    .trg_valid_i               (bound_trg_valid_o_6),
    .trg_ready_o               (bound_trg_ready_i_6),
    .trg_data_o                (bound_trg_data_i_6),
    .trg_valid_o               (bound_trg_valid_i_6),
    .trg_ready_i               (bound_trg_ready_o_6),
    .itp_data_i                (bound_itp_data_o_6),
    .itp_valid_i               (bound_itp_valid_o_6),
    .itp_ready_o               (bound_itp_ready_i_6),
    .itp_data_o                (bound_itp_data_i_6),
    .itp_valid_o               (bound_itp_valid_i_6),
    .itp_ready_i               (bound_itp_ready_o_6)
);

bound_link bl7(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_7),
    .trg_valid_i               (bound_trg_valid_o_7),
    .trg_ready_o               (bound_trg_ready_i_7),
    .trg_data_o                (bound_trg_data_i_7),
    .trg_valid_o               (bound_trg_valid_i_7),
    .trg_ready_i               (bound_trg_ready_o_7),
    .itp_data_i                (bound_itp_data_o_7),
    .itp_valid_i               (bound_itp_valid_o_7),
    .itp_ready_o               (bound_itp_ready_i_7),
    .itp_data_o                (bound_itp_data_i_7),
    .itp_valid_o               (bound_itp_valid_i_7),
    .itp_ready_i               (bound_itp_ready_o_7)
);

bound_link bl8(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_8),
    .trg_valid_i               (bound_trg_valid_o_8),
    .trg_ready_o               (bound_trg_ready_i_8),
    .trg_data_o                (bound_trg_data_i_8),
    .trg_valid_o               (bound_trg_valid_i_8),
    .trg_ready_i               (bound_trg_ready_o_8),
    .itp_data_i                (bound_itp_data_o_8),
    .itp_valid_i               (bound_itp_valid_o_8),
    .itp_ready_o               (bound_itp_ready_i_8),
    .itp_data_o                (bound_itp_data_i_8),
    .itp_valid_o               (bound_itp_valid_i_8),
    .itp_ready_i               (bound_itp_ready_o_8)
);

bound_link bl9(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_9),
    .trg_valid_i               (bound_trg_valid_o_9),
    .trg_ready_o               (bound_trg_ready_i_9),
    .trg_data_o                (bound_trg_data_i_9),
    .trg_valid_o               (bound_trg_valid_i_9),
    .trg_ready_i               (bound_trg_ready_o_9),
    .itp_data_i                (bound_itp_data_o_9),
    .itp_valid_i               (bound_itp_valid_o_9),
    .itp_ready_o               (bound_itp_ready_i_9),
    .itp_data_o                (bound_itp_data_i_9),
    .itp_valid_o               (bound_itp_valid_i_9),
    .itp_ready_i               (bound_itp_ready_o_9)
);

bound_link bl10(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_10),
    .trg_valid_i               (bound_trg_valid_o_10),
    .trg_ready_o               (bound_trg_ready_i_10),
    .trg_data_o                (bound_trg_data_i_10),
    .trg_valid_o               (bound_trg_valid_i_10),
    .trg_ready_i               (bound_trg_ready_o_10),
    .itp_data_i                (bound_itp_data_o_10),
    .itp_valid_i               (bound_itp_valid_o_10),
    .itp_ready_o               (bound_itp_ready_i_10),
    .itp_data_o                (bound_itp_data_i_10),
    .itp_valid_o               (bound_itp_valid_i_10),
    .itp_ready_i               (bound_itp_ready_o_10)
);

bound_link bl11(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_11),
    .trg_valid_i               (bound_trg_valid_o_11),
    .trg_ready_o               (bound_trg_ready_i_11),
    .trg_data_o                (bound_trg_data_i_11),
    .trg_valid_o               (bound_trg_valid_i_11),
    .trg_ready_i               (bound_trg_ready_o_11),
    .itp_data_i                (bound_itp_data_o_11),
    .itp_valid_i               (bound_itp_valid_o_11),
    .itp_ready_o               (bound_itp_ready_i_11),
    .itp_data_o                (bound_itp_data_i_11),
    .itp_valid_o               (bound_itp_valid_i_11),
    .itp_ready_i               (bound_itp_ready_o_11)
);

bound_link bl12(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_12),
    .trg_valid_i               (bound_trg_valid_o_12),
    .trg_ready_o               (bound_trg_ready_i_12),
    .trg_data_o                (bound_trg_data_i_12),
    .trg_valid_o               (bound_trg_valid_i_12),
    .trg_ready_i               (bound_trg_ready_o_12),
    .itp_data_i                (bound_itp_data_o_12),
    .itp_valid_i               (bound_itp_valid_o_12),
    .itp_ready_o               (bound_itp_ready_i_12),
    .itp_data_o                (bound_itp_data_i_12),
    .itp_valid_o               (bound_itp_valid_i_12),
    .itp_ready_i               (bound_itp_ready_o_12)
);

bound_link bl13(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_13),
    .trg_valid_i               (bound_trg_valid_o_13),
    .trg_ready_o               (bound_trg_ready_i_13),
    .trg_data_o                (bound_trg_data_i_13),
    .trg_valid_o               (bound_trg_valid_i_13),
    .trg_ready_i               (bound_trg_ready_o_13),
    .itp_data_i                (bound_itp_data_o_13),
    .itp_valid_i               (bound_itp_valid_o_13),
    .itp_ready_o               (bound_itp_ready_i_13),
    .itp_data_o                (bound_itp_data_i_13),
    .itp_valid_o               (bound_itp_valid_i_13),
    .itp_ready_i               (bound_itp_ready_o_13)
);

bound_link bl14(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_14),
    .trg_valid_i               (bound_trg_valid_o_14),
    .trg_ready_o               (bound_trg_ready_i_14),
    .trg_data_o                (bound_trg_data_i_14),
    .trg_valid_o               (bound_trg_valid_i_14),
    .trg_ready_i               (bound_trg_ready_o_14),
    .itp_data_i                (bound_itp_data_o_14),
    .itp_valid_i               (bound_itp_valid_o_14),
    .itp_ready_o               (bound_itp_ready_i_14),
    .itp_data_o                (bound_itp_data_i_14),
    .itp_valid_o               (bound_itp_valid_i_14),
    .itp_ready_i               (bound_itp_ready_o_14)
);

bound_link bl15(
    .clk                       (clk),
    .rstn                      (rstn),
    .trg_data_i                (bound_trg_data_o_15),
    .trg_valid_i               (bound_trg_valid_o_15),
    .trg_ready_o               (bound_trg_ready_i_15),
    .trg_data_o                (bound_trg_data_i_15),
    .trg_valid_o               (bound_trg_valid_i_15),
    .trg_ready_i               (bound_trg_ready_o_15),
    .itp_data_i                (bound_itp_data_o_15),
    .itp_valid_i               (bound_itp_valid_o_15),
    .itp_ready_o               (bound_itp_ready_i_15),
    .itp_data_o                (bound_itp_data_i_15),
    .itp_valid_o               (bound_itp_valid_i_15),
    .itp_ready_i               (bound_itp_ready_o_15)
);
endmodule
